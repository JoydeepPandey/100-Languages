// Hello World program in VERILOG
// Language: verilog
// File extension: .v

module hello;
    initial begin
        $display("Hello, World!");
        $finish;
    end
endmodule